library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity rom_and is
  Port (
    and_out : out std_logic_vector(3 downto 0);
    a : in std_logic_vector(3 downto 0);
    b : in std_logic_vector(3 downto 0) 
   );
end rom_and;

architecture Behavioral of rom_and is

--type rom is array (0 to 15) of std_logic_vector(1 downto 0 );
--signal memory : rom := ("00", "01", "10", "11", "01", "00", "11", "10", "10", "11", "00" , "01", "11", "10", "01", "00");
--signal addr : std_logic_vector(3 downto 0);


type rom_and is array (0 to 255) of std_logic_vector(3 downto 0 );
constant memory : rom_and := ("0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0000","0001", --17
"0000","0001","0000","0001","0000","0001","0000","0001","0000","0001","0000","0001","0000","0001","0000","0000","0010","0010","0000","0000","0010","0010","0000",
"0000","0010","0010","0000","0000","0010","0010","0000","0001","0010","0011","0000","0001","0010","0011","0000","0001","0010","0011","0000","0001","0010","0011",
"0000","0000","0000","0000","0100","0100","0100","0100","0000","0000","0000","0000","0100","0100","0100","0100","0000","0001","0000","0001","0100","0101","0100",
"0101","0000","0001","0000","0001","0100","0101","0100","0101","0000","0000","0010","0010","0100","0100","0110","0110","0000","0000","0010","0010","0100","0100",
"0110","0110","0000","0001","0010","0011","0100","0101","0110","0111","0000","0001","0010","0011","0100","0101","0110","0111","0000","0000","0000","0000","0000",
"0000","0000","0000","1000","1000","1000","1000","1000","1000","1000","1000","0000","0001","0000","0001","0000","0001","0000","0001","1000","1001","1000","1001",
"1000","1001","1000","1001","0000","0000","0010","0010","0000","0000","0010","0010","1000","1000","1010","1010","1000","1000","1010","1010","0000","0001","0010",
"0011","0000","0001","0010","0011","1000","1001","1010","1011","1000","1001","1010","1011","0000","0000","0000","0000","0100","0100","0100","0100","1000","1000",
"1000","1000","1100","1100","1100","1100","0000","0001","0000","0001","0100","0101","0100","0101","1000","1001","1000","1001","1100","1101","1100","1101","0000",
"0000","0010","0010","0100","0100","0110","0110","1000","1000","1010","1010","1100","1100","1110","1110","0000","0001","0010","0011","0100","0101","0110","0111",
"1000","1001","1010","1011","1100","1101","1110","1111");

signal addr : std_logic_vector(7 downto 0);
begin

addr <= a & b;
and_out <= memory(to_integer(unsigned(addr)));


end Behavioral;
