library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity rom_sigmoid is
  Port (
    sigmoid_out : out std_logic_vector(7 downto 0);
    a : in std_logic_vector(3 downto 0);
    b : in std_logic_vector(3 downto 0)
   );
end rom_sigmoid;

architecture Behavioral of rom_sigmoid is
--rom elements are not correct in this code.
type rom_sigmoid is array (0 to 255) of std_logic_vector(7 downto 0 );
constant memory : rom_sigmoid := ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000","00010000", --17
"00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00000000","00100000","00100000","00000000","00000000","00100000","00100000","00000000",

"00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00000000","00100000","00100000","00000000","00000000","00100000","00100000","00000000",

"00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00000000","00100000","00100000","00000000","00000000","00100000","00100000","00000000",

"00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00000000","00100000","00100000","00000000","00000000","00100000","00100000","00000000",

"00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00000000","00100000","00100000","00000000","00000000","00100000","00100000","00000000",

"00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00000000","00100000","00100000","00000000","00000000","00100000","00100000","00000000",

"00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00000000","00100000","00100000","00000000","00000000","00100000","00100000","00000000",

"00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00000000","00100000","00100000","00000000","00000000","00100000","00100000","00000000",

"00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00000000","00100000","00100000","00000000","00000000","00100000","00100000","00000000",
 
"00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00010000","00000000","00000000","00100000","00100000","00000000","00000000","00100000","00100000","00000000",

"10000000","10010000","10100000","10110000","11000000","11010000","11100000","11110000");

--"0000","0010","0010","0000","0000","0010","0010","0000","0001","0010","0011","0000","0001","0010","0011","0000","0001","0010","0011","0000","0001","0010","0011",
--"0000","0000","0000","0000","0100","0100","0100","0100","0000","0000","0000","0000","0100","0100","0100","0100","0000","0001","0000","0001","0100","0101","0100",
--"0101","0000","0001","0000","0001","0100","0101","0100","0101","0000","0000","0010","0010","0100","0100","0110","0110","0000","0000","0010","0010","0100","0100",
--"0110","0110","0000","0001","0010","0011","0100","0101","0110","0111","0000","0001","0010","0011","0100","0101","0110","0111","0000","0000","0000","0000","0000",
--"0000","0000","0000","1000","1000","1000","1000","1000","1000","1000","1000","0000","0001","0000","0001","0000","0001","0000","0001","1000","1001","1000","1001",
--"1000","1001","1000","1001","0000","0000","0010","0010","0000","0000","0010","0010","1000","1000","1010","1010","1000","1000","1010","1010","0000","0001","0010",
--"0011","0000","0001","0010","0011","1000","1001","1010","1011","1000","1001","1010","1011","0000","0000","0000","0000","0100","0100","0100","0100","1000","1000",
--"1000","1000","1100","1100","1100","1100","0000","0001","0000","0001","0100","0101","0100","0101","1000","1001","1000","1001","1100","1101","1100","1101","0000",
--"0000","0010","0010","0100","0100","0110","0110","1000","1000","1010","1010","1100","1100","1110","1110","0000","0001","0010","0011","0100","0101","0110","0111",
--"1000","1001","1010","1011","1100","1101","1110","1111");

signal addr : std_logic_vector(7 downto 0);
begin

addr <= a & b;
sigmoid_out <= memory(to_integer(unsigned(addr)));


end Behavioral;